module gf180mcu_bt_ip__logo;
endmodule
