module gf180mcu_bt_ip__tap;
endmodule
